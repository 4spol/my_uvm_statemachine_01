interface my_if (input  clk,input  rst_n);
	logic  vaild;
	logic  data;
endinterface

/*___________input interface____________*/
