interface my_ifo (input  clk,input  rst_n) ;
	logic en;
	logic [2:0]cnt;
	logic vaild;
endinterface

/*_________output interface______________*/